
package async_fifo_pkg;

`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "defines.sv"

`include "async_fifo_write_sequence_item.sv"
`include "async_fifo_read_sequence_item.sv"

`include "async_fifo_write_seq.sv"
`include "async_fifo_read_seq.sv"

`include "write_sequencer.sv"
`include "read_sequencer.sv"


`include "write_driver.sv"
`include "read_driver.sv"

`include "write_monitor.sv"
`include "read_monitor.sv"

`include "write_agent.sv"
`include "read_agent.sv"

`include "subscriber.sv"
`include "scoreboard.sv"

`include "virtual_sequencer.sv"

`include "environment.sv"
`include "virtual_sequence.sv"

`include "test.sv"


endpackage
